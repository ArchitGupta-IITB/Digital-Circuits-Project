library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity mem_blk is
	port(
		MEM_ADD: in std_logic_vector(15 downto 0);
		MEM_DATA_IN: in std_logic_vector(15 downto 0);
		--MEM_RD: in std_logic;
		MEM_WR: in std_logic;
		MEM_DATA_OUT: out std_logic_vector(15 downto 0)
	);
end entity mem_blk;

architecture mem_blk_bhv of mem_blk is
	--signals corresponding to 16-bit contents of 2^16 memory addresses need to be defined here
	type mem_vector is array (127 downto 0) of std_logic_vector(15 downto 0);
	signal MEM: mem_vector;
	signal MEM_DATA_TEMP: std_logic_vector(15 downto 0);
	signal index: integer;
	
begin
	index<=to_integer(unsigned(MEM_ADD));
	write_proc: process(index, MEM_WR, MEM_DATA_IN, MEM_ADD)
	begin
		--writing at negative edge in accordance with standard set in RF
			if(MEM_WR = '1') then
				MEM(to_integer(unsigned(MEM_ADD))) <= MEM_DATA_IN;
				--if statements need to be added for the other addresses
			end if;
		
	end process;
	
	read_proc: process(index, MEM_ADD)
	begin
		--if(clk'event and clk = '0') then
		--	if(MEM_RD = '1') then
				MEM_DATA_OUT <= MEM(to_integer(unsigned(MEM_ADD)));
				--if statements need to be added for the other addresses
			--end if;
		--end if;
	end process;
end architecture mem_blk_bhv;
		

 