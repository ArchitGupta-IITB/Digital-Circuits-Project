library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
<<<<<<< HEAD
=======

>>>>>>> 1c49dd2750449ff81e9fca3bce98eee2cac071c7
entity mem_blk is
	port(
		MEM_ADD: in std_logic_vector(15 downto 0);
		MEM_DATA_IN: in std_logic_vector(15 downto 0);
		MEM_RD: in std_logic;
		MEM_WR: in std_logic;
		clk: in std_logic;
		MEM_DATA_OUT: out std_logic_vector(15 downto 0)
	);
end entity mem_blk;

architecture mem_blk_bhv of mem_blk is
	--signals corresponding to 16-bit contents of 2^16 memory addresses need to be defined here
<<<<<<< HEAD
	signal MEM0: std_logic_vector(65535 downto 0);
=======
	type mem_vector is array (65535 downto 0) of std_logic_vector(15 downto 0);
	signal MEM: mem_vector;
>>>>>>> 1c49dd2750449ff81e9fca3bce98eee2cac071c7
	signal MEM_DATA_TEMP: std_logic_vector(15 downto 0);
	signal index: integer;
	
begin
	index<=to_integer(unsigned(MEM_ADD));
	write_proc: process(index, MEM_WR, clk)
	begin
		if(clk'event and clk = '0') then --writing at negative edge in accordance with standard set in RF
			if(MEM_WR = '1') then
<<<<<<< HEAD
				--index<=to_integer(unsigned(MEM_ADD));
				--if(MEM_ADD = "0000000000000000") then
					MEM0(index+15 downto index) <= MEM_DATA_IN;
				--end if;
=======
				MEM(to_integer(unsigned(MEM_ADD))) <= MEM_DATA_IN;
>>>>>>> 1c49dd2750449ff81e9fca3bce98eee2cac071c7
				--if statements need to be added for the other addresses
			end if;
		end if;
	end process;
	
	read_proc: process(index, MEM_RD, clk)
	begin
		if(clk'event and clk = '0') then
			if(MEM_RD = '1') then
<<<<<<< HEAD
				--if(MEM_ADD = "0000000000000000") then
					MEM_DATA_TEMP <= MEM0(index+15 downto index);
				--end if;
=======
				MEM_DATA_OUT <= MEM(to_integer(unsigned(MEM_ADD)));
>>>>>>> 1c49dd2750449ff81e9fca3bce98eee2cac071c7
				--if statements need to be added for the other addresses
			end if;
		end if;
	end process;
end architecture mem_blk_bhv;
		

 