library ieee;
use ieee.std_logic_1164.all;


entity fsm is
port(reset,clock: in std_logic);
end fsm;

architecture bhv of fsm is
---------------Define state type here-----------------------------
type state is (s1, s2, s3, s4, s5, s6, s7, s8, s9, s10, s11, s12, s13,
                s14, s15, s16, s17, s18, s19, s20, s21, s22 ); -- Fill other states here
---------------Define signals of state type-----------------------

component ALUA_MUX is 
port(
    S_ALU_A : in std_logic;
    RF_DA_OUT1 : in std_logic_vector(15 downto 0);
    T1 : in std_logic_vector(15 downto 0);ALUA_IN : out std_logic_vector(15 downto 0));
end component ALUA_MUX;

component ALUB_MUX is 
    port(
        --select signal
        S_ALU_B : in std_logic_vector(1 downto 0);

        -- input data
        PLUS1 : in std_logic_vector(15 downto 0);
        T2: in std_logic_vector(15 downto 0);
        SE16_6: in std_logic_vector(15 downto 0);
        SE16_9: in std_logic_vector(15 downto 0);
        --output data
        ALUB_IN : out std_logic_vector(15 downto 0)
    );
end component ALUB_MUX;

component ALU is
    port (
        ALU_A: in std_logic_vector(15 downto 0);
        ALU_B: in std_logic_vector(15 downto 0);
		alu_control: in std_logic_vector(1 downto 0);
        ALU_C: out std_logic_vector(15 downto 0);
		C: out std_logic;
		Z: out std_logic
    ) ;
end component ALU;

component IR_MUX is 
    port(
        --select signal
        S_IR : in std_logic;

        -- input data
        MEM_DATA_IR: in std_logic_vector(15 downto 0);
        LU_IR  : in std_logic_vector(15 downto 0);

        --output data
        IR_IN : out std_logic_vector(15 downto 0)

    );
end component IR_MUX;

component IR is
	port(
		IR_IN: in std_logic_vector(15 downto 0);
		IR_EN: in std_logic;
		IR_53: out std_logic_vector(2 downto 0);
		IR_86: out std_logic_vector(2 downto 0);
		IR_119: out std_logic_vector(2 downto 0);
		IR_50: out std_logic_vector(5 downto 0);
		IR_70: out std_logic_vector(7 downto 0);
		IR_80: out std_logic_vector(8 downto 0)
	);
end component IR;

component MEM_DATA_MUX is 
    port(
        --select signal
        S_MEM_DATA : in std_logic;

        -- input data
        RF_DA_IN  : in std_logic_vector(15 downto 0);
        RF_DA_OUT1: in std_logic_vector(15 downto 0);

        --output data
        MEM_DATA_IN : out std_logic_vector(15 downto 0)

    );
end component MEM_DATA_MUX;

component MEM_ADD_MUX is 
    port(
        --select signal
        S_MEM_ADD : in std_logic_vector(1 downto 0);

        -- input data
        RF_DA_OUT1 : in std_logic_vector(15 downto 0);
        T1: in std_logic_vector(15 downto 0);
        RF_DA_OUT2 : in std_logic_vector(15 downto 0);

        --output data
        MEM_ADD_IN : out std_logic_vector(15 downto 0)

    );
end component MEM_ADD_MUX;

component mem_blk is
	port(
		MEM_ADD: in std_logic_vector(15 downto 0);
		MEM_DATA_IN: in std_logic_vector(15 downto 0);
		MEM_RD: in std_logic;
		MEM_WR: in std_logic;
		clk: in std_logic;
		MEM_DATA_OUT: out std_logic_vector(15 downto 0)
	);
end component mem_blk;

component RF is 
    port(
        --to store the register number for each address
        RF_AD_OUT1 : in std_logic_vector(2 downto 0);
        RF_AD_OUT2 : in std_logic_vector(2 downto 0);
        RF_AD_IN : in std_logic_vector(2 downto 0);
        RF_reset: in std_logic;
        -- input data
        RF_DA_IN : in std_logic_vector(15 downto 0);

        RF_WR : in std_logic;
        --output data
        RF_DA_OUT1 : out std_logic_vector(15 downto 0);
        RF_DA_OUT2 : out std_logic_vector(15 downto 0)
    );
end component RF;

component RF_AD_OUT1_MUX is 
    port(
        --select signal
        S_RF_AD_OUT1 : in std_logic_vector(1 downto 0);

        -- input data
        IR86: in std_logic_vector(2 downto 0);
        IR119  : in std_logic_vector(2 downto 0);
        PEN_O : in std_logic_vector(2 downto 0);
        --output data
        RF_AD_OUT1 : out std_logic_vector(2 downto 0)

    );
end component RF_AD_OUT1_MUX;

component RF_AD_IN_MUX is 
    port(
        --select signal
        S_RF_AD_IN : in std_logic_vector(2 downto 0);

        -- input data
        IR53: in std_logic_vector(2 downto 0);
        IR86: in std_logic_vector(2 downto 0);
        IR119  : in std_logic_vector(2 downto 0);
        PEN_O : in std_logic_vector(2 downto 0);
        --output data
        RF_AD_IN : out std_logic_vector(2 downto 0)

    );
end component RF_AD_IN_MUX;


component RF_DA_IN_MUX is 
    port(
        --select signal
        S_RF_DA_IN : in std_logic_vector(1 downto 0);

        -- input data
        ALU_C : in std_logic_vector(15 downto 0);
        T1 : in std_logic_vector(15 downto 0);
        MEM_DATA: in std_logic_vector(15 downto 0);
        RF_DA_OUT1: in std_logic_vector(15 downto 0); 
        --output data
        RF_DA_IN : out std_logic_vector(15 downto 0)

    );
end component RF_DA_IN_MUX;


component T1_MUX is 
    port(
        --select signal
        S_T1 : in std_logic_vector(1 downto 0);

        -- input data
        RF_DA_OUT1_T1 : in std_logic_vector(15 downto 0);
        ALUC_T1: in std_logic_vector(15 downto 0);
        SE16_6_T1  : in std_logic_vector(15 downto 0);

        --output data
        T1_IN : out std_logic_vector(15 downto 0)

    );
end component T1_MUX;

component T2_MUX is 
    port(
        --select signal
        S_T2 : in std_logic;

        -- input data
        RF_DA_OUT2 : in std_logic_vector(15 downto 0);
        SE16_6  : in std_logic_vector(15 downto 0);

        --output data
        T2_IN : out std_logic_vector(15 downto 0)

    );
end component T2_MUX;


signal state_present,state_next: state:=s1;
signal S_ALU_A, S_IR, S_T2, S_MEM_DATA, C, Z, RF_WR,IR_EN,MEM_RD,MEM_WR,RF_reset,clk: std_logic;
signal S_ALU_B, S_ALU, S_RF_AD_OUT1, S_RF_DA_IN, S_T1, S_MEM_ADD, alu_control: std_logic_vector(1 downto 0);
signal S_RF_AD_IN,RF_AD_OUT1,RF_AD_OUT2,RF_AD_IN, IR_53,IR_86,IR_119,PEN_O: std_logic_vector(2 downto 0);
signal ALUA_IN,ALUB_IN, ALU_C, RF_DA_OUT1,RF_DA_OUT2,RF_DA_IN,T1,T2, SE16_6, SE16_9, IR_R, MEM_DATA_OUT,MEM_DATA_IN, LU_OUT,MEM_ADD_IN : std_logic_vector(15 downto 0);
signal PLUS1: std_logic_vector(15 downto 0);
signal IR_50: std_logic_vector(5 downto 0);
signal IR_70: std_logic_vector(7 downto 0);
signal IR_80: std_logic_vector(8 downto 0);
signal opcode: std_logic_vector(3 downto 0);

begin
ALU_A: ALUA_MUX port map(S_ALU_A,RF_DA_OUT1,T1,ALUA_IN);
ALU_B: ALUB_MUX port map(S_ALU_B, PLUS1,T2,SE16_6,SE16_9,ALUB_IN);
ALU_P: ALU port map(ALUA_IN, ALUB_IN,alu_control, ALU_C, C, Z);
IR_M: IR_MUX port map(S_IR, MEM_DATA_OUT,LU_OUT,IR_R);
IR_D: IR port map(IR_R,IR_EN,IR_53,IR_86,IR_119,IR_50,IR_70,IR_80);
RF1: RF port map(RF_AD_OUT1,RF_AD_OUT2,RF_AD_IN,RF_reset,RF_DA_IN,RF_WR,RF_DA_OUT1,RF_DA_OUT2);
RF_AD_IN_C: RF_AD_IN_MUX port map(S_RF_AD_IN,IR_53,IR_86,IR_119,PEN_O,RF_AD_IN);
RF_OUT1: RF_AD_OUT1_MUX port map(S_RF_AD_OUT1,IR_86,IR_119,PEN_O,RF_AD_OUT1);
RF_DA_IN_C: RF_DA_IN_MUX port map(S_RF_DA_IN,ALU_C,T1,MEM_DATA_OUT,RF_DA_OUT1,RF_DA_IN);
MEM_AD: MEM_ADD_MUX port map(S_MEM_ADD,RF_DA_OUT1,T1,RF_DA_OUT2,MEM_ADD_IN);
MEM_DA: MEM_DATA_MUX port map(S_MEM_DATA,RF_DA_IN,RF_DA_OUT1,MEM_DATA_IN);
MEM_BL: mem_blk port map(MEM_ADD_IN,MEM_DATA_IN,MEM_RD,MEM_WR,clk,MEM_DATA_OUT);
T1_M: T1_MUX port map(S_T1,RF_DA_OUT1,ALU_C,SE16_6,T1);
T2_M: T2_MUX port map(S_T2, RF_DA_OUT2,SE16_6,T2);
opcode<=IR_R(15 downto 12);
RF_AD_OUT2<=IR_119;

clock_proc:process(clock,reset)
    begin

        if(reset='1') then
        state_present<=s1;
        else
        if(clock='1' and clock' event) then
        state_present<=state_next;
        end if;
    end if;
end process;


state_transition_proc:process(state_present,opcode)
begin
case state_present is
    when s1=>
    S_RF_AD_OUT1 <= "00";
    S_IR<='0';
    S_RF_AD_IN<="000";
    S_RF_DA_IN<="00";
    S_MEM_ADD<= "00";
    S_IR<='0';
    if(opcode = "0000" or opcode = "0010" or opcode = "0001" or
        opcode = "0100" or opcode = "0101" or opcode = "1100") then-- Fill the code here
        state_next<=s2;
    elsif(opcode ="0011" ) then--FILL OTHER STATES HERE
        state_next<=s7;
    elsif(opcode = "1000") then
        state_next<=s12;
    elsif(opcode ="1001") then
        state_next<=s16;
    elsif(opcode = "0110") then
        state_next<=s18;
    elsif(opcode= "0111") then
        state_next<=s22;
    else
        state_next<=s1;
    end if;

    when s2=>
    S_RF_AD_OUT1<="01";
    S_T1<="00";
    if(opcode = "0000" or opcode = "0001") then
        state_next<=s3; -- Fill the code here
        S_T2<='0';
    elsif (opcode = "0100" or opcode = "0101") then
        state_next<=s3;
        S_T2<='1';
    elsif(opcode = "0010") then
        state_next<=s5;
        S_T2<='0';
    elsif(opcode = "1100") then
        state_next<=s11;
    else
        state_next<=s1;
    end if;
    when s3=>
    S_ALU_A<='1';
    S_ALU_B<="01";
    S_T1<="01";
    if(opcode = "0000") then
        state_next<=s4; 
    elsif(opcode = "0001") then
        state_next<=s6;
    elsif(opcode = "0100") then
        state_next<=s9;
    elsif(opcode = "0101") then
        state_next<=s10;
    else
        state_next<=s1;
    end if;
    when s4=>
        state_next<=s1;
        S_RF_AD_IN<="001"; 
        S_RF_DA_IN<="01";

    when s5=>
        state_next<=s4;
        S_ALU_A<='1';
        S_ALU_B<="01";
        S_T1<="01";

    when s6=>
        state_next<=s1;
        S_RF_AD_IN<="010";
        S_RF_DA_IN<="01";
    when s7=>
        state_next<=s8;
        S_T1<="10";    
    when s8=>
        state_next<=s1;
        S_RF_AD_IN<="011";
        S_RF_DA_IN<="01";

    when s9=>
        state_next<=s1;
        S_MEM_DATA<='0';
        S_MEM_ADD<="01";
        S_RF_DA_IN<="10";
        S_RF_AD_IN<="011";
    when s10=>
        state_next<=s1;
        S_RF_AD_OUT1<="10";
        S_MEM_ADD<="01";
        S_MEM_DATA<='1';

    when s11=>
        S_T1<="01";
        S_ALU_B<="01";
        S_ALU_A<='1';
        if( Z = '1') then
            state_next<=s12;
        else
            state_next<=s1;
        end if;
    
    when s12=>
        S_ALU_A<='0';
        S_ALU_B<="00";
        S_RF_AD_OUT1<="00";
        S_RF_AD_IN<="000";
        S_RF_DA_IN<= "00";

        if(opcode = "1100") then
            state_next<=s13;
        elsif(opcode = "1000") then
            state_next<=s14;
        else
            state_next<=s1;
        end if;

    when s13=>
        state_next<=s1;
        S_ALU_A<= '0';
        S_ALU_B<="10";
        S_RF_AD_OUT1<="00";
        S_RF_AD_IN<="000";
        S_RF_DA_IN<="00";

    when s14=>
        state_next<=s15;

        S_RF_AD_OUT1<="00";    
        S_RF_AD_IN<="011";
        S_RF_DA_IN<="11";
    
    when s15=>
        state_next<=s1;

        S_ALU_A<='0';
        S_ALU_B<="11";
        S_RF_AD_OUT1<="00";
        S_RF_AD_IN<="000";
        S_RF_DA_IN<="00";

    when s16=>
        state_next<=s17;
        S_ALU_A<='0';
        S_ALU_B<="00";
        S_RF_AD_OUT1<="00";
        S_RF_AD_IN<="011";
        S_RF_DA_IN<="00";

    when s17=>
        state_next<=s1;
        S_RF_AD_OUT1<="01";
        S_RF_AD_IN<="000";
        S_RF_DA_IN<="11";
    when s18=>
            
        if( Z= '0') then
            state_next<=s19;
        else
            state_next<=s1;
        end if;
    
    when s19=>  
        state_next<=s20;
        S_RF_AD_OUT1<="10";
        S_RF_AD_IN<="100";
        S_RF_DA_IN<="10";
        S_T1<="00";
        S_MEM_ADD<="00";
        S_MEM_DATA<='0';
        S_IR<='1';
    when s20=>
        S_IR<='0';
        S_RF_DA_IN<="00";
        S_RF_AD_IN<="011";
        S_ALU_A<='1';
        S_ALU_B<="00";
        if(opcode = "0110") then
            state_next<=s18;
        elsif(opcode = "0111") then
            state_next<=s22;
        else
            state_next<=s1;
        end if;
    
    when s22=>
           
        if(Z = '0') then
            state_next<=s21;
        else
            state_next<=s1;
        end if;

    when s21=>
        state_next<=s20;
        S_MEM_DATA<='1';
        S_MEM_ADD<="10";
        S_RF_AD_OUT1<="11";
        S_IR<='1';
    when others=>
        state_next<=s1;
    
end case;
end process;

-------------------------
---------Fill rest of the code here---------

end bhv;
